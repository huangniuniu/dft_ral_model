`ifndef _RAL_DEFINE_SVH
`define _RAL_DEFINE_SVH

//------------------------------------------------------------------------------
//TDR definition

//==========add by hcai1 for mtap1149 TDR begin=================//
`define IEEE_1149_WBYPASS_OPCODE           `IEEE_1149_IR_WIDTH'h00
`define IEEE_1149_WBYPASS_LENGTH            1
`define IEEE_1149_WBYPASS_RST_VALUE        `IEEE_1149_WBYPASS_LENGTH'h0
`define IEEE_1149_WBYPASS_ADDR             {`IEEE_1149_WBYPASS_OPCODE,`SIB_WIDTH'h0} 

`define IEEE_1149_PIPELINEMODE_OPCODE     `IEEE_1149_IR_WIDTH'h01
`define IEEE_1149_PIPELINEMODE_LENGTH      1
`define IEEE_1149_PIPELINEMODE_RST_VALUE   `IEEE_1149_PIPELINEMODE_LENGTH'h0
`define IEEE_1149_PIPELINEMODE_ADDR        {`IEEE_1149_PIPELINEMODE_OPCODE,`SIB_WIDTH'h0} 

`define IEEE_1149_IDCODE_OPCODE           `IEEE_1149_IR_WIDTH'h02
`define IEEE_1149_IDCODE_LENGTH            32
`define IEEE_1149_IDCODE_RST_VALUE        `IEEE_1149_IDCODE_LENGTH'h3
`define IEEE_1149_IDCODE_ADDR             {`IEEE_1149_IDCODE_OPCODE,`SIB_WIDTH'h0}

`define IEEE_1149_MANID_OPCODE           `IEEE_1149_IR_WIDTH'h1f
`define IEEE_1149_MANID_LENGTH            28
`define IEEE_1149_MANID_RST_VALUE        `IEEE_1149_MANID_LENGTH'h3
`define IEEE_1149_MANID_ADDR             {`IEEE_1149_MANID_OPCODE,`SIB_WIDTH'h0}

`define SOC_STAC_WBYPASS_OPCODE           `IEEE_1500_IR_WIDTH'h00
`define SOC_STAC_WBYPASS_LENGTH            1
`define SOC_STAC_WBYPASS_RST_VALUE        `SOC_STAC_WBYPASS_LENGTH'h0
`define SOC_STAC_WBYPASS_ADDR             {`SOC_STAC_WBYPASS_OPCODE,`SIB_WIDTH'h1} 

`define SOC_STAC_BYPASS_OPCODE           `IEEE_1500_IR_WIDTH'hff
`define SOC_STAC_BYPASS_LENGTH            1
`define SOC_STAC_BYPASS_RST_VALUE        `SOC_STAC_BYPASS_LENGTH'h0
`define SOC_STAC_BYPASS_ADDR             {`SOC_STAC_BYPASS_OPCODE,`SIB_WIDTH'h1}

`define SOC_STAC_MEMCFG_OPCODE           `IEEE_1500_IR_WIDTH'h76
`define SOC_STAC_MEMCFG_LENGTH            22
`define SOC_STAC_MEMCFG_RST_VALUE        `SOC_STAC_MEMCFG_LENGTH'h0
`define SOC_STAC_MEMCFG_ADDR             {`SOC_STAC_MEMCFG_OPCODE,`SIB_WIDTH'h1}

`define SOC_STAC_IOCTRL_OPCODE           `IEEE_1500_IR_WIDTH'h73
`define SOC_STAC_IOCTRL_LENGTH            14
`define SOC_STAC_IOCTRL_RST_VALUE        `SOC_STAC_IOCTRL_LENGTH'h0
`define SOC_STAC_IOCTRL_ADDR             {`SOC_STAC_IOCTRL_OPCODE,`SIB_WIDTH'h1}

//==========add by hcai1 for mtap1149 TDR end===================//


`define SCANCONFIG_OPCODE         `IEEE_1500_IR_WIDTH'h24
`define SCANCONFIG_LENGTH         14
`define SCANCONFIG_RST_VALUE      `SCANCONFIG_LENGTH'h6c
//`define SCANCONFIG_ADDR           {`SCANCONFIG_OPCODE,`SIB_WIDTH'b0010} 
`define SCANCONFIG_ADDR           `DFT_REG_ADDR_WIDTH'h242  

`define IDCODE_OPCODE         `IEEE_1500_IR_WIDTH'hfc
`define IDCODE_LENGTH         8
`define IDCODE_RST_VALUE      `IDCODE_LENGTH'h6c
`define IDCODE_ADDR           {`IDCODE_OPCODE,`SIB_WIDTH'b0101} 

`define BYPASS_OPCODE         `IEEE_1149_IR_WIDTH'hff
`define BYPASS_LENGTH         1
`define BYPASS_RST_VALUE      `BYPASS_LENGTH'h0
`define BYPASS_ADDR          {`BYPASS_OPCODE,`SIB_WIDTH'h0} 

`define P1687_OPCODE         `IEEE_1149_IR_WIDTH'h13
`define P1687_LENGTH         `LVL1SIB_WIDTH 
`define P1687_RST_VALUE      `P1687_LENGTH'h0
`define P1687_ADDR           {`P1687_OPCODE,`SIB_WIDTH'h0} 

`define SUB_CLIENT_SIB_OPCODE         `IEEE_1500_IR_WIDTH'h13
`define SUB_CLIENT_SIB_LENGTH         `LVL2SIB_WIDTH 
`define SUB_CLIENT_SIB_RST_VALUE      `SUB_CLIENT_SIB_LENGTH'h0
`define SUB_CLIENT_SIB_ADDR           {`SUB_CLIENT_SIB_OPCODE,`SIB_WIDTH'h1} 

`define P1687_QRYUPD_ONLY_OPCODE    `IEEE_1500_IR_WIDTH'h14

`define DUMMY_TDR_OPCODE         `IEEE_1149_IR_WIDTH'h3c
`define DUMMY_TDR_ADDR          {`DUMMY_TDR_OPCODE,`SIB_WIDTH'h0} 
`define DUMMY_TDR_LENGTH         350
`define DUMMY_TDR_FIELD1_WIDTH   100
`define DUMMY_TDR_FIELD1_RST_VALUE `DUMMY_TDR_FIELD1_WIDTH'hff
`define DUMMY_TDR_FIELD2_WIDTH   100
`define DUMMY_TDR_FIELD2_RST_VALUE `DUMMY_TDR_FIELD1_WIDTH'h55
`define DUMMY_TDR_FIELD3_WIDTH   150
`define DUMMY_TDR_FIELD3_RST_VALUE `DUMMY_TDR_FIELD1_WIDTH'haa

//------------------------------------------------------------------------------
//Master TAP ALTTAPEN
//------------------------------------------------------------------------------
`define MTAP_ALTTAPEN_OPCODE         `IEEE_1149_IR_WIDTH'h5
`define MTAP_ALTTAPEN_ADDR           {`MTAP_ALTTAPEN_OPCODE,`SIB_WIDTH'h0} 
`define MTAP_ALTTAPEN_LENGTH         4
`define MTAP_ALTTAPEN_RST_VALUE      0

//------------------------------------------------------------------------------
//GOPPHY_CRSEL Define
//------------------------------------------------------------------------------
`define GOPPHY_CRSEL_OPCODE                  `GOPPHY_IR_WIDTH'h31
`define GOPPHY_CRSEL_ADDR                    {`GOPPHY_CRSEL_OPCODE,`SIB_WIDTH'h0} 
`define GOPPHY_CRSEL_LENGTH                  18
`define GOPPHY_CRSEL_ADD_DATA_WIDTH          16
`define GOPPHY_CRSEL_ADD_DATA_RST_VALUE      `GOPPHY_CRSEL_ADD_DATA_WIDTH'h0 
`define GOPPHY_CRSEL_CMD_WIDTH               2
`define GOPPHY_CRSEL_CMD_RST_VALUE           `GOPPHY_CRSEL_ADD_DATA_WIDTH'h0 


//------------------------------------------------------------------------------
//SoC STAC ALTTAPEN
//------------------------------------------------------------------------------
`define SOC_STAC_ALTTAPEN_OPCODE                      `IEEE_1500_IR_WIDTH'h5
`define SOC_STAC_ALTTAPEN_ADDR                        {`SOC_STAC_ALTTAPEN_OPCODE,`SIB_WIDTH'h1} 
`define SOC_STAC_ALTTAPEN_LENGTH                      9 
`define SOC_STAC_ALTTAPEN_RST_VALUE                   0
`define SOC_STAC_ALTTAPEN_SOC_STAC_WIDTH              1 
`define SOC_STAC_ALTTAPEN_SOC_STAC_RST_VALUE          0 
`define SOC_STAC_ALTTAPEN_GOPPHYX2_STAC_WIDTH              1 
`define SOC_STAC_ALTTAPEN_GOPPHYX2_STAC_RST_VALUE          0 

//------------------------------------------------------------------------------
//LVL2 1687
//------------------------------------------------------------------------------
`define LVL2_P1687_OPCODE         `IEEE_1500_IR_WIDTH'h13
`define LVL2_P1687_LENGTH         `LVL2SIB_WIDTH 
`define LVL2_P1687_RST_VALUE      `LVL2_P1687_LENGTH'h0
`define LVL2_P1687_ADDR           {`LVL2_P1687_OPCODE,`SIB_WIDTH'1} 
//------------------------------------------------------------------------------
//SYSPLL_CFG_TDR Define
//------------------------------------------------------------------------------
`define SYSPLL1_CFG_OPCODE         `IEEE_1500_IR_WIDTH'h60
`define SYSPLL2_CFG_OPCODE         `IEEE_1500_IR_WIDTH'h61
`define SYSPLL_CFG_LENGTH         400
`define SYSPLL_CFG_RST_VALUE      `SYSPLL_CFG_LENGTH'h0
`define SYSPLL1_CFG_LENGTH         400
`define SYSPLL1_CFG_RST_VALUE      `SYSPLL1_CFG_LENGTH'h0
`define SYSPLL2_CFG_LENGTH         400
`define SYSPLL2_CFG_RST_VALUE      `SYSPLL2_CFG_LENGTH'h0
`define SYSPLL1_CFG_ADDR           {`SYSPLL1_CFG_OPCODE,`SIB_WIDTH'h1} 
//BOZO: SYSPLL2_CFG_OPCODE has not released thus far.
`define SYSPLL2_CFG_ADDR           {`SYSPLL2_CFG_OPCODE,`SIB_WIDTH'h1} 

//------------------------------------------------------------------------------
//DPLL1_CSRACCESS Define
//------------------------------------------------------------------------------
`define DPLL1_CSRACCESS_OPCODE         `IEEE_1500_IR_WIDTH'h62
`define DPLL1_CSRACCESS_LENGTH         51
`define DPLL1_CSRACCESS_RST_VALUE      `DPLL1_CSRACCESS_LENGTH'h0
`define DPLL1_CSRACCESS_ADDR           {`DPLL1_CSRACCESS_OPCODE,`SIB_WIDTH'b1} 
`define DPLL1_CSRACCESS_COMPLETE_RD_WR_WIDTH       1
`define DPLL1_CSRACCESS_COMPLETE_RD_WR_LSB         0
`define DPLL1_CSRACCESS_COMPLETE_RD_WR_RST_VALUE   `DPLL1_CSRACCESS_COMPLETE_RD_WR_WIDTH'h0
`define DPLL1_CSRACCESS_CFG_DATA_WIDTH       32
`define DPLL1_CSRACCESS_CFG_DATA_LSB         `DPLL1_CSRACCESS_COMPLETE_RD_WR_LSB+`DPLL1_CSRACCESS_COMPLETE_RD_WR_WIDTH
`define DPLL1_CSRACCESS_CFG_DATA_RST_VALUE   `DPLL1_CSRACCESS_COMPLETE_RD_WR_WIDTH'h0
`define DPLL1_CSRACCESS_CFG_ADDR_WIDTH       16
`define DPLL1_CSRACCESS_CFG_ADDR_LSB         `DPLL1_CSRACCESS_CFG_DATA_LSB+`DPLL1_CSRACCESS_CFG_DATA_WIDTH
`define DPLL1_CSRACCESS_CFG_ADDR_RST_VALUE   `DPLL1_CSRACCESS_CFG_ADDR_WIDTH'h0
`define DPLL1_CSRACCESS_EXECUTE_WIDTH       1
`define DPLL1_CSRACCESS_EXECUTE_LSB         `DPLL1_CSRACCESS_CFG_ADDR_LSB+`DPLL1_CSRACCESS_CFG_ADDR_WIDTH
`define DPLL1_CSRACCESS_EXECUTE_RST_VALUE   `DPLL1_CSRACCESS_EXECUTE_WIDTH'h0
`define DPLL1_CSRACCESS_CFG_PROTECTB_WIDTH       1
`define DPLL1_CSRACCESS_CFG_PROTECTB_LSB         `DPLL1_CSRACCESS_EXECUTE_LSB+`DPLL1_CSRACCESS_EXECUTE_WIDTH
`define DPLL1_CSRACCESS_CFG_PROTECTB_RST_VALUE   `DPLL1_CSRACCESS_CFG_PROTECTB_WIDTH'h0

//------------------------------------------------------------------------------
//TESTCONFIG_TDR Define
//------------------------------------------------------------------------------
`define TESTCONFIG_OPCODE         `IEEE_1500_IR_WIDTH'h67
`define TESTCONFIG_LENGTH         33
`define TESTCONFIG_RST_VALUE      `TESTCONFIG_LENGTH'h0
`define TESTCONFIG_ADDR           {`TESTCONFIG_OPCODE,`SIB_WIDTH'b1} 
`define TESTCONFIG_PLLBYPASSEN_WIDTH       1
`define TESTCONFIG_PLLBYPASSEN_LSB         0
`define TESTCONFIG_PLLBYPASSEN_RST_VALUE   `TESTCONFIG_PLLBYPASSEN_WIDTH'h0
`define TESTCONFIG_PFH_SCAN_SCANMODE_WIDTH       4
`define TESTCONFIG_PFH_SCAN_SCANMODE_LSB         `TESTCONFIG_PLLBYPASSEN_LSB+`TESTCONFIG_PLLBYPASSEN_WIDTH
`define TESTCONFIG_PFH_SCAN_SCANMODE_RST_VALUE   `TESTCONFIG_PFH_SCAN_SCANMODE_WIDTH'h0
`define TESTCONFIG_TILE_TESTMODE1_WIDTH       1
`define TESTCONFIG_TILE_TESTMODE1_LSB         `TESTCONFIG_PFH_SCAN_SCANMODE_LSB+`TESTCONFIG_PFH_SCAN_SCANMODE_WIDTH
`define TESTCONFIG_TILE_TESTMODE1_RST_VALUE   `TESTCONFIG_TILE_TESTMODE1_WIDTH'h0
`define TESTCONFIG_TILE_TESTMODE2_WIDTH       1
`define TESTCONFIG_TILE_TESTMODE2_LSB         `TESTCONFIG_TILE_TESTMODE1_LSB+`TESTCONFIG_TILE_TESTMODE1_WIDTH
`define TESTCONFIG_TILE_TESTMODE2_RST_VALUE   `TESTCONFIG_TILE_TESTMODE2_WIDTH'h0
`define TESTCONFIG_TILE_TESTMODE3_WIDTH       1
`define TESTCONFIG_TILE_TESTMODE3_LSB         `TESTCONFIG_TILE_TESTMODE2_LSB+`TESTCONFIG_TILE_TESTMODE2_WIDTH
`define TESTCONFIG_TILE_TESTMODE3_RST_VALUE   `TESTCONFIG_TILE_TESTMODE3_WIDTH'h0
`define TESTCONFIG_OCC_TESTMODE_WIDTH       1
`define TESTCONFIG_OCC_TESTMODE_LSB         `TESTCONFIG_TILE_TESTMODE3_LSB+`TESTCONFIG_TILE_TESTMODE3_WIDTH
`define TESTCONFIG_OCC_TESTMODE_RST_VALUE   `TESTCONFIG_OCC_TESTMODE_WIDTH'h0
`define TESTCONFIG_SCANMODE_WIDTH       1
`define TESTCONFIG_SCANMODE_LSB         `TESTCONFIG_OCC_TESTMODE_LSB+`TESTCONFIG_OCC_TESTMODE_WIDTH
`define TESTCONFIG_SCANMODE_RST_VALUE   `TESTCONFIG_SCANMODE_WIDTH'h0
`define TESTCONFIG_TILE_SEL_WIDTH       18
`define TESTCONFIG_TILE_SEL_LSB         `TESTCONFIG_SCANMODE_LSB+`TESTCONFIG_SCANMODE_WIDTH
`define TESTCONFIG_TILE_SEL_RST_VALUE   `TESTCONFIG_TILE_SEL_WIDTH'h0
`define TESTCONFIG_RESERVE_WIDTH       5
`define TESTCONFIG_RESERVE_LSB         `TESTCONFIG_TILE_SEL_LSB+`TESTCONFIG_TILE_SEL_WIDTH
`define TESTCONFIG_RESERVE_RST_VALUE   `TESTCONFIG_RESERVE_WIDTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_TESTMODE Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_TESTMODE_OPCODE         `IEEE_1500_IR_WIDTH'h46
`define GOPPHY_DFT_GASKET_2_LANECONFIG_TESTMODE_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_TESTMODE_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_TESTMODE_LENGTH         30
`define GOPPHY_DFT_GASKET_2_LANECONFIG_TESTMODE_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_TESTMODE_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_ALTTAP_EN Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_ALTTAP_EN_OPCODE             `IEEE_1500_IR_WIDTH'h05
`define GOPPHY_DFT_GASKET_2_ALTTAP_EN_ADDR               {`GOPPHY_DFT_GASKET_2_ALTTAP_EN_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_ALTTAP_EN_LENGTH             2
`define GOPPHY_DFT_GASKET_2_ALTTAP_EN_SIPC0_WIDTH        1
`define GOPPHY_DFT_GASKET_2_ALTTAP_EN_SIPC0_RST_VALUE    0 
`define GOPPHY_DFT_GASKET_2_ALTTAP_EN_ENABLE_WIDTH       1
`define GOPPHY_DFT_GASKET_2_ALTTAP_EN_ENABLE_RST_VALUE   0 

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_TESTMODE Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_TESTMODE_OPCODE         `IEEE_1500_IR_WIDTH'h46
`define GOPPHY_DFT_GASKET_4_LANECONFIG_TESTMODE_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_TESTMODE_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_TESTMODE_LENGTH         390
`define GOPPHY_DFT_GASKET_4_LANECONFIG_TESTMODE_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_TESTMODE_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_ALTTAP_EN Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_ALTTAP_EN_OPCODE             `IEEE_1500_IR_WIDTH'h05
`define GOPPHY_DFT_GASKET_4_ALTTAP_EN_ADDR               {`GOPPHY_DFT_GASKET_4_ALTTAP_EN_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_ALTTAP_EN_LENGTH             2
`define GOPPHY_DFT_GASKET_4_ALTTAP_EN_SIPC0_WIDTH        1
`define GOPPHY_DFT_GASKET_4_ALTTAP_EN_SIPC0_RST_VALUE    0 
`define GOPPHY_DFT_GASKET_4_ALTTAP_EN_ENABLE_WIDTH       1
`define GOPPHY_DFT_GASKET_4_ALTTAP_EN_ENABLE_RST_VALUE   0 

//gaowei begin add macro define for GOP*2 TDRs and GOP*4 TDRs
//below is for GOP2
//GOPPHY_DFT_GASKET_2_LANECONFIG_SCANCONFIG Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_SCANCONFIG_OPCODE         `IEEE_1500_IR_WIDTH'h09
`define GOPPHY_DFT_GASKET_2_LANECONFIG_SCANCONFIG_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_SCANCONFIG_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_SCANCONFIG_LENGTH         18
`define GOPPHY_DFT_GASKET_2_LANECONFIG_SCANCONFIG_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_SCANCONFIG_LENGTH'hb0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_CLOCK_SELECT Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLOCK_SELECT_OPCODE         `IEEE_1500_IR_WIDTH'h4c
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLOCK_SELECT_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_CLOCK_SELECT_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLOCK_SELECT_LENGTH         2
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLOCK_SELECT_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_CLOCK_SELECT_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_CLK_OBSERVE Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLK_OBSERVE_OPCODE         `IEEE_1500_IR_WIDTH'h4d
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLK_OBSERVE_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_CLK_OBSERVE_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLK_OBSERVE_LENGTH         28
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CLK_OBSERVE_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_CLK_OBSERVE_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_ANALOG_OBS_EN Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ANALOG_OBS_EN_OPCODE         `IEEE_1500_IR_WIDTH'h4e
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ANALOG_OBS_EN_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_ANALOG_OBS_EN_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ANALOG_OBS_EN_LENGTH         3
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ANALOG_OBS_EN_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_ANALOG_OBS_EN_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_CHANNEL_BYPASS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CHANNEL_BYPASS_OPCODE         `IEEE_1500_IR_WIDTH'h4f
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CHANNEL_BYPASS_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_CHANNEL_BYPASS_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CHANNEL_BYPASS_LENGTH         4
`define GOPPHY_DFT_GASKET_2_LANECONFIG_CHANNEL_BYPASS_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_CHANNEL_BYPASS_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_COUNTER Define 
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_COUNTER_OPCODE         `IEEE_1500_IR_WIDTH'h50
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_COUNTER_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_COUNTER_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_COUNTER_LENGTH         8
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_COUNTER_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_COUNTER_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_ROSEN Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_ROSEN_OPCODE         `IEEE_1500_IR_WIDTH'h51
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_ROSEN_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_ROSEN_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_ROSEN_LENGTH         1
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_ROSEN_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_CNTL_ROSEN_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_SETUP Define 
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_SETUP_OPCODE         `IEEE_1500_IR_WIDTH'h52
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_SETUP_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_SETUP_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_SETUP_LENGTH         9
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_SETUP_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_SETUP_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_STATUS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_STATUS_OPCODE         `IEEE_1500_IR_WIDTH'h53
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_STATUS_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_STATUS_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_STATUS_LENGTH         30
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_STATUS_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_ROS_STATUS_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_OPCODE         `IEEE_1500_IR_WIDTH'h56
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_LENGTH         97
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_STATUS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_STATUS_OPCODE         `IEEE_1500_IR_WIDTH'h57
`define GOPPHY_DFT_GASKET_2_LANECONFIG_STATUS_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_STATUS_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_STATUS_LENGTH         25//gaowei 26 in doc
`define GOPPHY_DFT_GASKET_2_LANECONFIG_STATUS_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_STATUS_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_BSR_DEBUG Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_BSR_DEBUG_OPCODE         `IEEE_1500_IR_WIDTH'h47
`define GOPPHY_DFT_GASKET_2_LANECONFIG_BSR_DEBUG_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_BSR_DEBUG_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_BSR_DEBUG_LENGTH         10
`define GOPPHY_DFT_GASKET_2_LANECONFIG_BSR_DEBUG_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_BSR_DEBUG_LENGTH'h0

//------------------------------------------------------------------------------

//GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_OPCODE         `IEEE_1500_IR_WIDTH'h56
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_LENGTH         97
`define GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_MPLL_CONTROL_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_OPCODE         `IEEE_1500_IR_WIDTH'h49
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_LENGTH         69
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RX Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RX_OPCODE         `IEEE_1500_IR_WIDTH'h4a
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RX_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RX_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RX_LENGTH         33
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RX_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_RX_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_TX Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_TX_OPCODE         `IEEE_1500_IR_WIDTH'h4b
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_TX_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_TX_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_TX_LENGTH         41
`define GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_TX_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_LOOPBACK_TX_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_CTRL Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_CTRL_OPCODE         `IEEE_1500_IR_WIDTH'h58
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_CTRL_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_CTRL_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_CTRL_LENGTH         41
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_CTRL_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_CTRL_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_OBS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_OBS_OPCODE         `IEEE_1500_IR_WIDTH'h59
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_OBS_ADDR           {`GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_OBS_OPCODE,`SIB_WIDTH'h3} 
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_OBS_LENGTH         17
`define GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_OBS_RST_VALUE      `GOPPHY_DFT_GASKET_2_LANECONFIG_ISOLATION_CHAIN_OBS_LENGTH'h0
//finish GOP2


//below is for GOP4
//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_SCANCONFIG Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_SCANCONFIG_OPCODE         `IEEE_1500_IR_WIDTH'h09
`define GOPPHY_DFT_GASKET_4_LANECONFIG_SCANCONFIG_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_SCANCONFIG_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_SCANCONFIG_LENGTH         18
`define GOPPHY_DFT_GASKET_4_LANECONFIG_SCANCONFIG_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_SCANCONFIG_LENGTH'hb0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_BSR_DEBUG Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_BSR_DEBUG_OPCODE         `IEEE_1500_IR_WIDTH'h47
`define GOPPHY_DFT_GASKET_4_LANECONFIG_BSR_DEBUG_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_BSR_DEBUG_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_BSR_DEBUG_LENGTH         10
`define GOPPHY_DFT_GASKET_4_LANECONFIG_BSR_DEBUG_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_BSR_DEBUG_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_OPCODE         `IEEE_1500_IR_WIDTH'h49//gaowei 39 in doc
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_LENGTH         121
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_TX Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_TX_OPCODE         `IEEE_1500_IR_WIDTH'h4b
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_TX_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_TX_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_TX_LENGTH         41
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_TX_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_TX_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RX Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RX_OPCODE         `IEEE_1500_IR_WIDTH'h4a
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RX_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RX_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RX_LENGTH         33
`define GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RX_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_LOOPBACK_RX_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_COUNTER Define 
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_COUNTER_OPCODE         `IEEE_1500_IR_WIDTH'h50
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_COUNTER_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_COUNTER_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_COUNTER_LENGTH         8
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_COUNTER_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_COUNTER_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_ROSEN Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_ROSEN_OPCODE         `IEEE_1500_IR_WIDTH'h51
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_ROSEN_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_ROSEN_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_ROSEN_LENGTH         1
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_ROSEN_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_CNTL_ROSEN_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_SETUP Define 
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_SETUP_OPCODE         `IEEE_1500_IR_WIDTH'h52
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_SETUP_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_SETUP_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_SETUP_LENGTH         9
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_SETUP_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_SETUP_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_STATUS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_STATUS_OPCODE         `IEEE_1500_IR_WIDTH'h53
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_STATUS_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_STATUS_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_STATUS_LENGTH         30
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_STATUS_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_ROS_STATUS_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_MPLL_CONTROL Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_MPLL_CONTROL_OPCODE         `IEEE_1500_IR_WIDTH'h56
`define GOPPHY_DFT_GASKET_4_LANECONFIG_MPLL_CONTROL_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_MPLL_CONTROL_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_MPLL_CONTROL_LENGTH         97
`define GOPPHY_DFT_GASKET_4_LANECONFIG_MPLL_CONTROL_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_MPLL_CONTROL_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_STATUS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_STATUS_OPCODE         `IEEE_1500_IR_WIDTH'h57
`define GOPPHY_DFT_GASKET_4_LANECONFIG_STATUS_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_STATUS_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_STATUS_LENGTH         25//gaowei 26 in doc
`define GOPPHY_DFT_GASKET_4_LANECONFIG_STATUS_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_STATUS_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_CTRL Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_CTRL_OPCODE         `IEEE_1500_IR_WIDTH'h58
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_CTRL_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_CTRL_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_CTRL_LENGTH         41
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_CTRL_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_CTRL_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_OBS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_OBS_OPCODE         `IEEE_1500_IR_WIDTH'h59
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_OBS_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_OBS_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_OBS_LENGTH         17
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_OBS_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_ISOLATION_CHAIN_OBS_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_CLOCK_SELECT Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLOCK_SELECT_OPCODE         `IEEE_1500_IR_WIDTH'h4c
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLOCK_SELECT_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_CLOCK_SELECT_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLOCK_SELECT_LENGTH         2
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLOCK_SELECT_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_CLOCK_SELECT_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_CLK_OBSERVE Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLK_OBSERVE_OPCODE         `IEEE_1500_IR_WIDTH'h4d
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLK_OBSERVE_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_CLK_OBSERVE_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLK_OBSERVE_LENGTH         42
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CLK_OBSERVE_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_CLK_OBSERVE_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_CHANNEL_BYPASS Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CHANNEL_BYPASS_OPCODE         `IEEE_1500_IR_WIDTH'h4f
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CHANNEL_BYPASS_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_CHANNEL_BYPASS_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CHANNEL_BYPASS_LENGTH         5
`define GOPPHY_DFT_GASKET_4_LANECONFIG_CHANNEL_BYPASS_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_CHANNEL_BYPASS_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ANALOG_OBS_EN Define
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ANALOG_OBS_EN_OPCODE         `IEEE_1500_IR_WIDTH'h4e
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ANALOG_OBS_EN_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_ANALOG_OBS_EN_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ANALOG_OBS_EN_LENGTH         3
`define GOPPHY_DFT_GASKET_4_LANECONFIG_ANALOG_OBS_EN_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_ANALOG_OBS_EN_LENGTH'h0

//------------------------------------------------------------------------------
//GOPPHY_DFT_GASKET_4_LANECONFIG_ Define  for 00/ff I-bass
//------------------------------------------------------------------------------
`define GOPPHY_DFT_GASKET_4_LANECONFIG_WS_BYPASS_OPCODE         `IEEE_1500_IR_WIDTH'h00
`define GOPPHY_DFT_GASKET_4_LANECONFIG_WS_BYPASS_ADDR           {`GOPPHY_DFT_GASKET_4_LANECONFIG_WS_BYPASS_OPCODE,`SIB_WIDTH'h5} 
`define GOPPHY_DFT_GASKET_4_LANECONFIG_WS_BYPASS_LENGTH         1
`define GOPPHY_DFT_GASKET_4_LANECONFIG_WS_BYPASS_RST_VALUE      `GOPPHY_DFT_GASKET_4_LANECONFIG_WS_BYPASS_LENGTH'h0

//gaowei end


//------------------------------------------------------------------------------
//TMDPPHY_1_CFGACCESS Define
//------------------------------------------------------------------------------
`define TMDPPHY_1_CFGACCESS_OPCODE         `IEEE_1500_IR_WIDTH'h41
`define TMDPPHY_1_CFGACCESS_ADDR           {`TMDPPHY_1_CFGACCESS_OPCODE,`SIB_WIDTH'h9} 
`define TMDPPHY_1_CFGACCESS_LENGTH         50
`define TMDPPHY_1_CFGACCESS_RST_VALUE      `TMDPPHY_1_CFGACCESS_LENGTH'h0

//------------------------------------------------------------------------------
//TMDPPHY_1_SCANCONFIG Define
//------------------------------------------------------------------------------
`define TMDPPHY_1_SCANCONFIG_OPCODE         `IEEE_1500_IR_WIDTH'h9
`define TMDPPHY_1_SCANCONFIG_ADDR           {`TMDPPHY_1_SCANCONFIG_OPCODE,`SIB_WIDTH'h9} 
`define TMDPPHY_1_SCANCONFIG_LENGTH         17
`define TMDPPHY_1_SCANCONFIG_RST_VALUE      `TMDPPHY_1_SCANCONFIG_LENGTH'h0


`define PLLCFG_OPCODE         `IEEE_1149_IR_WIDTH'h60
`define PLLCFG_LENGTH         400
`define PLLCFG_RST_VALUE      `PLLCFG_LENGTH'h0
`define PLLCFG_ADDR           {`PLLCFG_OPCODE,`SIB_WIDTH'h1} 

//Child STC 1687 OPCODE
`define P1687A_OPCODE         `IEEE_1149_IR_WIDTH'h13
`define MANID_OPCODE          `IEEE_1149_IR_WIDTH'h1F


//FUSE_OVERRIDE TDR Define
`define FUSE_OVERRIDE_OPCODE         `IEEE_1500_IR_WIDTH'h74
`define FUSE_OVERRIDE_LENGTH         512
`define FUSE_OVERRIDE_RST_VALUE      `FUSE_OVERRIDE_LENGTH'h0
`define FUSE_OVERRIDE_ADDR           {`FUSE_OVERRIDE_OPCODE,`SIB_WIDTH'h1} 
`define FUSE_OVERRIDE_FIELD1_WIDTH   512
`define FUSE_OVERRIDE_FIELD1_RST_VALUE `FUSE_OVERRIDE_FIELD1_WIDTH'h0

//SPTAP_JPC_WIR TDR Define
`define SPTAP_JPC_WIR_OPCODE         3'b001
//`define SPTAP_JPC_WIR_LENGTH         6
//`define SPTAP_JPC_WIR_RST_VALUE      `SPTAP_JPC_WIR_LENGTH'h0
//`define SPTAP_JPC_WIR_ADDR           {`SPTAP_JPC_WIR_OPCODE,`SIB_WIDTH'h0} 
//SPTAP_JPC_WDR TDR Define
`define SPTAP_JPC_WDR_OPCODE         3'b010
//`define SPTAP_JPC_WDR_LENGTH         512
//`define SPTAP_JPC_WDR_RST_VALUE      `SPTAP_JPC_WDR_LENGTH'h0
//`define SPTAP_JPC_WDR_ADDR           {`SPTAP_JPC_WDR_OPCODE,`SIB_WIDTH'h0} 
//SPTAP_SMS_WIR TDR Define
`define SPTAP_SMS_WIR_OPCODE         3'b011
//`define SPTAP_SMS_WIR_LENGTH         6
//`define SPTAP_SMS_WIR_RST_VALUE      `SPTAP_SMS_WIR_LENGTH'h0
//`define SPTAP_SMS_WIR_ADDR           {`SPTAP_SMS_WIR_OPCODE,`SIB_WIDTH'h0} 
//SPTAP_SMS_WDR TDR Define
`define SPTAP_SMS_WDR_OPCODE         3'b100
//`define SPTAP_SMS_WDR_LENGTH         32
//`define SPTAP_SMS_WDR_RST_VALUE      `SPTAP_SMS_WDR_LENGTH'h0
//`define SPTAP_SMS_WDR_ADDR           {`SPTAP_SMS_WDR_OPCODE,`SIB_WIDTH'h0} 
//SPTAP BYPASS TDR Define
`define SPTAP_BYPASS_OPCODE    3'b111
`define SPTAP_BYPASS_LENGTH    1
`define SPTAP_BYPASS_RST_VALUE `SPTAP_BYPASS_LENGTH'h0
`define SPTAP_BYPASS_ADDR      {`SPTAP_BYPASS_OPCODE,`SIB_WIDTH'h0} 

//JPC_WIR TDR Define
`define JPC_WIR_OPCODE         `IEEE_1500_IR_WIDTH'h6d
//`define JPC_WIR_LENGTH         6
//`define JPC_WIR_RST_VALUE      `JPC_WIR_LENGTH'h0
//`define JPC_WIR_ADDR           {`JPC_WIR_OPCODE,`SIB_WIDTH'h1} 
//JPC_WDR TDR Define
`define JPC_WDR_OPCODE         `IEEE_1500_IR_WIDTH'h6e
//`define JPC_WDR_LENGTH         512
//`define JPC_WDR_RST_VALUE      `JPC_WDR_LENGTH'h0
//`define JPC_WDR_ADDR           {`JPC_WDR_OPCODE,`SIB_WIDTH'h1} 
//SMS_WIR TDR Define
`define SMS_WIR_OPCODE         `IEEE_1500_IR_WIDTH'h6f
//`define SMS_WIR_LENGTH         6
//`define SMS_WIR_RST_VALUE      `SMS_WIR_LENGTH'h0
//`define SMS_WIR_ADDR           {`SMS_WIR_OPCODE,`SIB_WIDTH'h1} 
//SMS_WDR TDR Define
`define SMS_WDR_OPCODE         `IEEE_1500_IR_WIDTH'h70
//`define SMS_WDR_LENGTH         32
//`define SMS_WDR_RST_VALUE      `SMS_WDR_LENGTH'h0
//`define SMS_WDR_ADDR           {`SMS_WDR_OPCODE,`SIB_WIDTH'h1} 

//SMS_STATUS TDR Define
`define SMS_STATUS_OPCODE         `IEEE_1500_IR_WIDTH'h71
`define SMS_STATUS_LENGTH         51
`define SMS_STATUS_RST_VALUE      `SMS_STATUS_LENGTH'h0
`define SMS_STATUS_ADDR           {`SMS_STATUS_OPCODE,`SIB_WIDTH'h1} 
//SMS_CONFIG TDR Define
`define SMS_CONFIG_OPCODE         `IEEE_1500_IR_WIDTH'h72
`define SMS_CONFIG_LENGTH         61
`define SMS_CONFIG_RST_VALUE      `SMS_CONFIG_LENGTH'h0
`define SMS_CONFIG_ADDR           {`SMS_CONFIG_OPCODE,`SIB_WIDTH'h1}

//gaowei add define for lvds
//LVDS_SERDES TDR Define
`define LVDS_SERDES_OPCODE        `IEEE_1500_IR_WIDTH'h77
`define LVDS_SERDES_LENGTH        14
`define LVDS_SERDES_RST_VALUE     `LVDS_SERDES_LENGTH'h0
`define LVDS_SERDES_ADDR          {`LVDS_SERDES_OPCODE,`SIB_WIDTH'h1} 
//LVDS_APB TDR Define
`define LVDS_APB_OPCODE          `IEEE_1500_IR_WIDTH'h78
`define LVDS_APB_LENGTH          21
`define LVDS_APB_RST_VALUE       `LVDS_APB_LENGTH'h0
`define LVDS_APB_ADDR            {`LVDS_APB_OPCODE,`SIB_WIDTH'h1}



//SPTAP JPC TDR define
`define SPTAP_JPC_SMS_SEL_OPCODE         `SMS_IR_WIDTH'h21
`define SPTAP_JPC_SMS_SEL_LENGTH         5
`define SPTAP_JPC_SMS_SEL_RST_VALUE      `SPTAP_JPC_SMS_SEL_LENGTH'h0
`define SPTAP_JPC_SMS_SEL_ADDR           {`SPTAP_JPC_SMS_SEL_OPCODE,`SPTAP_JPC_TDR} 

`define SPTAP_JPC_UDR_SEL_OPCODE         `SMS_IR_WIDTH'h35
`define SPTAP_JPC_UDR_SEL_LENGTH         512
`define SPTAP_JPC_UDR_SEL_RST_VALUE      `SPTAP_JPC_UDR_SEL_LENGTH'h0
`define SPTAP_JPC_UDR_SEL_ADDR           {`SPTAP_JPC_UDR_SEL_OPCODE,`SPTAP_JPC_TDR} 

//SPTAP SMS TDR define
`define SPTAP_SMS_TBOX_SEL_OPCODE         `SMS_IR_WIDTH'h2
`define SPTAP_SMS_TBOX_SEL_LENGTH         151
`define SPTAP_SMS_TBOX_SEL_RST_VALUE      `SPTAP_SMS_TBOX_SEL_LENGTH'h0
`define SPTAP_SMS_TBOX_SEL_ADDR           {`SPTAP_SMS_TBOX_SEL_OPCODE,`SPTAP_SMS_TDR} 

//JPC TDR define
`define JPC_SMS_SEL_OPCODE         `SMS_IR_WIDTH'h21
`define JPC_SMS_SEL_LENGTH         5
`define JPC_SMS_SEL_RST_VALUE      `JPC_SMS_SEL_LENGTH'h0
`define JPC_SMS_SEL_ADDR           {`JPC_SMS_SEL_OPCODE,`MTAP_JPC_TDR} 

`define JPC_BR_SEL_OPCODE         `SMS_IR_WIDTH'h2a
`define JPC_BR_SEL_LENGTH         6
`define JPC_BR_SEL_RST_VALUE      `JPC_BR_SEL_LENGTH'h0
`define JPC_BR_SEL_ADDR           {`JPC_BR_SEL_OPCODE,`MTAP_JPC_TDR} 

`define JPC_UDR_SEL_OPCODE         `SMS_IR_WIDTH'h35
`define JPC_UDR_SEL_LENGTH         512
`define JPC_UDR_SEL_RST_VALUE      `JPC_UDR_SEL_LENGTH'h0
`define JPC_UDR_SEL_ADDR           {`JPC_UDR_SEL_OPCODE,`MTAP_JPC_TDR} 

`define JPC_UDR_LOAD_OPCODE         `SMS_IR_WIDTH'h34
`define JPC_UDR_LOAD_LENGTH         6
`define JPC_UDR_LOAD_RST_VALUE      `JPC_UDR_LOAD_LENGTH'h0
`define JPC_UDR_LOAD_ADDR           {`JPC_UDR_LOAD_OPCODE,`MTAP_JPC_TDR} 

`define JPC_PGMR_SEL_OPCODE         `SMS_IR_WIDTH'h28
`define JPC_PGMR_SEL_LENGTH         12
`define JPC_PGMR_SEL_RST_VALUE      `JPC_PGMR_SEL_LENGTH'h0
`define JPC_PGMR_SEL_ADDR           {`JPC_PGMR_SEL_OPCODE,`MTAP_JPC_TDR} 

`define JPC_UDR_PROGRAM_OPCODE         `SMS_IR_WIDTH'h37
`define JPC_UDR_PROGRAM_LENGTH         6
`define JPC_UDR_PROGRAM_RST_VALUE      `JPC_UDR_PROGRAM_LENGTH'h0
`define JPC_UDR_PROGRAM_ADDR           {`JPC_UDR_PROGRAM_OPCODE,`MTAP_JPC_TDR} 

`define JPC_UDR_COMPARE_OPCODE         `SMS_IR_WIDTH'h36
`define JPC_UDR_COMPARE_LENGTH         6
`define JPC_UDR_COMPARE_RST_VALUE      `JPC_UDR_COMPARE_LENGTH'h0
`define JPC_UDR_COMPARE_ADDR           {`JPC_UDR_COMPARE_OPCODE,`MTAP_JPC_TDR} 

`define JPC_RBOX_RST_OPCODE         `SMS_IR_WIDTH'h24
`define JPC_RBOX_RST_LENGTH         6
`define JPC_RBOX_RST_RST_VALUE      `JPC_RBOX_RST_LENGTH'h0
`define JPC_RBOX_RST_ADDR           {`JPC_RBOX_RST_OPCODE,`MTAP_JPC_TDR} 

`define JPC_RBOX_SEL_OPCODE         `SMS_IR_WIDTH'h25
`define JPC_RBOX_SEL_LENGTH         512
`define JPC_RBOX_SEL_RST_VALUE      `JPC_RBOX_SEL_LENGTH'h0
`define JPC_RBOX_SEL_ADDR           {`JPC_RBOX_SEL_OPCODE,`MTAP_JPC_TDR} 

`define JPC_RBOX_PROGRAM_OPCODE         `SMS_IR_WIDTH'h27
`define JPC_RBOX_PROGRAM_LENGTH         6
`define JPC_RBOX_PROGRAM_RST_VALUE      `JPC_RBOX_PROGRAM_LENGTH'h0
`define JPC_RBOX_PROGRAM_ADDR           {`JPC_RBOX_PROGRAM_OPCODE,`MTAP_JPC_TDR} 

`define JPC_RBOX_COMPARE_OPCODE         `SMS_IR_WIDTH'h26
`define JPC_RBOX_COMPARE_LENGTH         6
`define JPC_RBOX_COMPARE_RST_VALUE      `JPC_RBOX_COMPARE_LENGTH'h0
`define JPC_RBOX_COMPARE_ADDR           {`JPC_RBOX_COMPARE_OPCODE,`MTAP_JPC_TDR} 

`define JPC_STATUS_SEL_OPCODE         `SMS_IR_WIDTH'h09
`define JPC_STATUS_SEL_LENGTH         6
`define JPC_STATUS_SEL_RST_VALUE      `JPC_STATUS_SEL_LENGTH'h0
`define JPC_STATUS_SEL_ADDR           {`JPC_STATUS_SEL_OPCODE,`MTAP_JPC_TDR} 

//SMS TDR define
`define SMS_TBOX_SEL_OPCODE         `SMS_IR_WIDTH'h2
`define SMS_TBOX_SEL_LENGTH         151
`define SMS_TBOX_SEL_RST_VALUE      `SMS_TBOX_SEL_LENGTH'h0
`define SMS_TBOX_SEL_ADDR           {`SMS_TBOX_SEL_OPCODE,`MTAP_SMS_TDR}

//GDDR5 IOCTRL define
`define GDDR5_IOCTRL_OPCODE        `IEEE_1500_IR_WIDTH'h73
`define GDDR5_IOCTRL_LENGTH        14
`define GDDR5_IOCTRL_RST_VALUE     `GDDR5_IOCTRL_LENGTH'h0
`define GDDR5_IOCTRL_ADDR          {`GDDR5_IOCTRL_OPCODE,`SIB_WIDTH'h1}
`endif
