`include "../top/ral_define.svh"
`include "../top/dft_reg.svh"
`include "../top/dft_reg_map.svh"
`include "../top/dft_reg_block.svh"
`include "../top/ral_class.sv"
