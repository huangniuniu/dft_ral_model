`ifndef _ASSIGN_SYSTEMPLL_DFT_SV
`define _ASSIGN_SYSTEMPLL_DFT_SV

    `define SPLL_PATH DUT.systempll_dft0

    assign  DUT.RefClk_p = pll_if.gen_spll_refclk_k;
    assign  DUT.RefClk_n =~pll_if.gen_spll_refclk_k;

    assign  pll_if.BP_ANALOG=                             `SPLL_PATH.BP_ANALOG;
    assign  `SPLL_PATH.gen_spll_alt_nctl=                 pll_if.gen_spll_alt_nctl;
    assign  `SPLL_PATH.gen_spll_alt_nctl_en=              pll_if.gen_spll_alt_nctl_en;
    assign  `SPLL_PATH.gen_spll_anaobs_sel=               pll_if.gen_spll_anaobs_sel;
    assign  `SPLL_PATH.gen_spll_bleeder_ac=               pll_if.gen_spll_bleeder_ac;
    assign  `SPLL_PATH.gen_spll_bleeder_en=               pll_if.gen_spll_bleeder_en;
    assign  `SPLL_PATH.gen_spll_bypass_freq_lock=         pll_if.gen_spll_bypass_freq_lock;
    assign  `SPLL_PATH.gen_spll_cfg_update_req=           pll_if.gen_spll_cfg_update_req;
    assign  `SPLL_PATH.gen_spll_clear_sticky_lock=        pll_if.gen_spll_clear_sticky_lock;
    assign  `SPLL_PATH.gen_spll_clk_nctl_sel=             pll_if.gen_spll_clk_nctl_sel;
    assign  `SPLL_PATH.gen_spll_clk_tdc_sel=              pll_if.gen_spll_clk_tdc_sel;
    assign  `SPLL_PATH.gen_spll_coarse_tdc_dis=           pll_if.gen_spll_coarse_tdc_dis;
    assign  `SPLL_PATH.gen_spll_dc_scan=                  pll_if.gen_spll_dc_scan;
    assign  `SPLL_PATH.gen_spll_dclk8_sel=                pll_if.gen_spll_dclk8_sel;
    assign  `SPLL_PATH.gen_spll_dco_cfg=                  pll_if.gen_spll_dco_cfg;
    assign  `SPLL_PATH.gen_spll_dft_capture=              pll_if.gen_spll_dft_capture;
    assign  `SPLL_PATH.gen_spll_dft_sel=                  pll_if.gen_spll_dft_sel;
    assign  `SPLL_PATH.gen_spll_digobs_div=               pll_if.gen_spll_digobs_div;
    assign  `SPLL_PATH.gen_spll_digobs_sel=               pll_if.gen_spll_digobs_sel;
    assign  `SPLL_PATH.gen_spll_digobs_trig_div=          pll_if.gen_spll_digobs_trig_div;
    assign  `SPLL_PATH.gen_spll_digobs_trig_sel=          pll_if.gen_spll_digobs_trig_sel;
    assign  `SPLL_PATH.gen_spll_divider_reset_refclk=     pll_if.gen_spll_divider_reset_refclk;
    assign  `SPLL_PATH.gen_spll_dpll_cfg_1=               pll_if.gen_spll_dpll_cfg_1;
    assign  `SPLL_PATH.gen_spll_dpll_cfg_2=               pll_if.gen_spll_dpll_cfg_2;
    assign  `SPLL_PATH.gen_spll_dpll_cfg_3=               pll_if.gen_spll_dpll_cfg_3;
    assign  `SPLL_PATH.gen_spll_duty_cycle_adj=           pll_if.gen_spll_duty_cycle_adj;
    assign  `SPLL_PATH.gen_spll_fb_slip_dis=              pll_if.gen_spll_fb_slip_dis;
    assign  `SPLL_PATH.gen_spll_fbclk_track_refclk=       pll_if.gen_spll_fbclk_track_refclk;
    assign  `SPLL_PATH.gen_spll_fbdiv_mask_en=            pll_if.gen_spll_fbdiv_mask_en;
    assign  `SPLL_PATH.gen_spll_fcw0_frac=                pll_if.gen_spll_fcw0_frac;
    assign  `SPLL_PATH.gen_spll_fcw0_int=                 pll_if.gen_spll_fcw0_int;
    assign  `SPLL_PATH.gen_spll_fcw1_frac=                pll_if.gen_spll_fcw1_frac;
    assign  `SPLL_PATH.gen_spll_fcw1_int=                 pll_if.gen_spll_fcw1_int;
    assign  `SPLL_PATH.gen_spll_fcw_denom=                pll_if.gen_spll_fcw_denom;
    assign  `SPLL_PATH.gen_spll_fcw_sel=                  pll_if.gen_spll_fcw_sel;
    assign  `SPLL_PATH.gen_spll_fcw_slew_frac=            pll_if.gen_spll_fcw_slew_frac;
    assign  `SPLL_PATH.gen_spll_fine_tdc_dis=             pll_if.gen_spll_fine_tdc_dis;
    assign  `SPLL_PATH.gen_spll_fracn_en=                 pll_if.gen_spll_fracn_en;
    assign  `SPLL_PATH.gen_spll_freq_jump_en=             pll_if.gen_spll_freq_jump_en;
    assign  `SPLL_PATH.gen_spll_gi_coarse_exp=            pll_if.gen_spll_gi_coarse_exp;
    assign  `SPLL_PATH.gen_spll_gi_coarse_mant=           pll_if.gen_spll_gi_coarse_mant;
    assign  `SPLL_PATH.gen_spll_gp_coarse_exp=            pll_if.gen_spll_gp_coarse_exp;
    assign  `SPLL_PATH.gen_spll_gp_coarse_mant=           pll_if.gen_spll_gp_coarse_mant;
    assign  `SPLL_PATH.gen_spll_is_1p2=                   pll_if.gen_spll_is_1p2;
    assign  `SPLL_PATH.gen_spll_iso_vddout_on_vddin=      pll_if.gen_spll_iso_vddout_on_vddin;
    assign  `SPLL_PATH.gen_spll_kdco_cal_dis=             pll_if.gen_spll_kdco_cal_dis;
    assign  `SPLL_PATH.gen_spll_kdco_incr_cal_dis=        pll_if.gen_spll_kdco_incr_cal_dis;
    assign  `SPLL_PATH.gen_spll_kdco_ratio=               pll_if.gen_spll_kdco_ratio;
    assign  `SPLL_PATH.gen_spll_lock_det_dis=             pll_if.gen_spll_lock_det_dis;
    assign  `SPLL_PATH.gen_spll_lock_det_tdc_steps=       pll_if.gen_spll_lock_det_tdc_steps;
    assign  `SPLL_PATH.gen_spll_lock_timer=               pll_if.gen_spll_lock_timer;
    assign  `SPLL_PATH.gen_spll_meas_win_sel=             pll_if.gen_spll_meas_win_sel;
    assign  `SPLL_PATH.gen_spll_misc_fuse_ctrl=           pll_if.gen_spll_misc_fuse_ctrl;
    assign  `SPLL_PATH.gen_spll_nctl_adj_dis=             pll_if.gen_spll_nctl_adj_dis;
    assign  `SPLL_PATH.gen_spll_nctl_coarse_frac_res=     pll_if.gen_spll_nctl_coarse_frac_res;
    assign  `SPLL_PATH.gen_spll_nctl_coarse_res=          pll_if.gen_spll_nctl_coarse_res;
    assign  `SPLL_PATH.gen_spll_nctl_coarse_step_dis=     pll_if.gen_spll_nctl_coarse_step_dis;
    assign  `SPLL_PATH.gen_spll_nctl_sig_del_dis=         pll_if.gen_spll_nctl_sig_del_dis;
    assign  `SPLL_PATH.gen_spll_pa_pll_test=              pll_if.gen_spll_pa_pll_test;
    assign  `SPLL_PATH.gen_spll_phase_jump_trig=          pll_if.gen_spll_phase_jump_trig;
    assign  `SPLL_PATH.gen_spll_phase_offset=             pll_if.gen_spll_phase_offset;
    assign  `SPLL_PATH.gen_spll_phy_analog_out=           pll_if.gen_spll_phy_analog_out;
    assign  `SPLL_PATH.gen_spll_pll_bypass=               pll_if.gen_spll_pll_bypass;
    assign  `SPLL_PATH.gen_spll_pll_bypass_clk=           pll_if.gen_spll_pll_bypass_clk;
    assign  `SPLL_PATH.gen_spll_pll_charz_ext_h=          pll_if.gen_spll_pll_charz_ext_h;
    assign  `SPLL_PATH.gen_spll_pll_charz_ext_l=          pll_if.gen_spll_pll_charz_ext_l;
    assign  `SPLL_PATH.gen_spll_pll_charz_sel=            pll_if.gen_spll_pll_charz_sel;
    assign  `SPLL_PATH.gen_spll_pll_en=                   pll_if.gen_spll_pll_en;
    assign  `SPLL_PATH.gen_spll_pll_test_en=              pll_if.gen_spll_pll_test_en;
    assign  `SPLL_PATH.gen_spll_pllout_req=               pll_if.gen_spll_pllout_req;
    assign  `SPLL_PATH.gen_spll_pllout_sel=               pll_if.gen_spll_pllout_sel;
    assign  `SPLL_PATH.gen_spll_pllout_state=             pll_if.gen_spll_pllout_state;
    assign  `SPLL_PATH.gen_spll_postdiv=                  pll_if.gen_spll_postdiv;
    assign  `SPLL_PATH.gen_spll_postdiv_pllout=           pll_if.gen_spll_postdiv_pllout;
    assign  `SPLL_PATH.gen_spll_postdiv_req=              pll_if.gen_spll_postdiv_req;
    assign  `SPLL_PATH.gen_spll_postdiv_sync_enable=      pll_if.gen_spll_postdiv_sync_enable;
    assign  `SPLL_PATH.gen_spll_prbs_en=                  pll_if.gen_spll_prbs_en;
    assign  `SPLL_PATH.gen_spll_pulse_mode=               pll_if.gen_spll_pulse_mode;
    assign  `SPLL_PATH.gen_spll_pwr_good=                 pll_if.gen_spll_pwr_good;
    assign  `SPLL_PATH.gen_spll_pwr_state=                pll_if.gen_spll_pwr_state;
    assign  `SPLL_PATH.gen_spll_pwrok_vddin=              pll_if.gen_spll_pwrok_vddin;
    assign  `SPLL_PATH.gen_spll_pwrok_vddout=             pll_if.gen_spll_pwrok_vddout;
    assign  `SPLL_PATH.gen_spll_refclk_bypass_vddout=     pll_if.gen_spll_refclk_bypass_vddout;
    assign  `SPLL_PATH.gen_spll_refclk_div=               pll_if.gen_spll_refclk_div;
    assign  `SPLL_PATH.gen_spll_refclk_gate_dis=          pll_if.gen_spll_refclk_gate_dis;
    //temp assign  `SPLL_PATH.gen_spll_refclk_k=                 pll_if.gen_spll_refclk_k;
    assign  `SPLL_PATH.gen_spll_refclk_rate=              pll_if.gen_spll_refclk_rate;
    assign  `SPLL_PATH.gen_spll_reg_obs_sel=              pll_if.gen_spll_reg_obs_sel;
    assign  `SPLL_PATH.gen_spll_reg_off_hi=               pll_if.gen_spll_reg_off_hi;
    assign  `SPLL_PATH.gen_spll_reg_off_lo=               pll_if.gen_spll_reg_off_lo;
    assign  `SPLL_PATH.gen_spll_reg_on_mode=              pll_if.gen_spll_reg_on_mode;
    assign  `SPLL_PATH.gen_spll_rlad_tap_sel=             pll_if.gen_spll_rlad_tap_sel;
    assign  `SPLL_PATH.gen_spll_scale_driver=             pll_if.gen_spll_scale_driver;
    assign  `SPLL_PATH.gen_spll_scan_clk=                 pll_if.gen_spll_scan_clk;
    assign  `SPLL_PATH.gen_spll_scan_in=                  pll_if.gen_spll_scan_in;
    assign  `SPLL_PATH.gen_spll_scan_shift_en=            pll_if.gen_spll_scan_shift_en;
    assign  `SPLL_PATH.gen_spll_sel_bump=                 pll_if.gen_spll_sel_bump;
    assign  `SPLL_PATH.gen_spll_sel_rladder_x=            pll_if.gen_spll_sel_rladder_x;
    assign  `SPLL_PATH.gen_spll_shrink_clk=               pll_if.gen_spll_shrink_clk;
    assign  `SPLL_PATH.gen_spll_shrink_mode=              pll_if.gen_spll_shrink_mode;
    assign  `SPLL_PATH.gen_spll_sig_del_patt_sel=         pll_if.gen_spll_sig_del_patt_sel;
    assign  `SPLL_PATH.gen_spll_ssc_en=                   pll_if.gen_spll_ssc_en;
    assign  `SPLL_PATH.gen_spll_stop_clk=                 pll_if.gen_spll_stop_clk;
    assign  `SPLL_PATH.gen_spll_stop_mode=                pll_if.gen_spll_stop_mode;
    assign  `SPLL_PATH.gen_spll_stop_mode_select=         pll_if.gen_spll_stop_mode_select;
    assign  `SPLL_PATH.gen_spll_syncbus_his_en=           pll_if.gen_spll_syncbus_his_en;
    assign  `SPLL_PATH.gen_spll_syncbus_in_refclk=        pll_if.gen_spll_syncbus_in_refclk;
    assign  `SPLL_PATH.gen_spll_tdc_cal_ctrl=             pll_if.gen_spll_tdc_cal_ctrl;
    assign  `SPLL_PATH.gen_spll_tdc_cal_en=               pll_if.gen_spll_tdc_cal_en;
    assign  `SPLL_PATH.gen_spll_tdc_clk_gate_en=          pll_if.gen_spll_tdc_clk_gate_en;
    assign  `SPLL_PATH.gen_spll_tdc_resolution=           pll_if.gen_spll_tdc_resolution;
    assign  `SPLL_PATH.gen_spll_trig_coarse_step=         pll_if.gen_spll_trig_coarse_step;
    assign  pll_if.spll_gen_dclk4_0=                      `SPLL_PATH.spll_gen_dclk4_0;
    assign  pll_if.spll_gen_dclk4_180=                    `SPLL_PATH.spll_gen_dclk4_180;
    assign  pll_if.spll_gen_dclk4_270=                    `SPLL_PATH.spll_gen_dclk4_270;
    assign  pll_if.spll_gen_dclk4_90=                     `SPLL_PATH.spll_gen_dclk4_90;
    assign  pll_if.spll_gen_dclk8_0=                      `SPLL_PATH.spll_gen_dclk8_0;
    assign  pll_if.spll_gen_dclk8_135=                    `SPLL_PATH.spll_gen_dclk8_135;
    assign  pll_if.spll_gen_dclk8_180=                    `SPLL_PATH.spll_gen_dclk8_180;
    assign  pll_if.spll_gen_dclk8_225=                    `SPLL_PATH.spll_gen_dclk8_225;
    assign  pll_if.spll_gen_dclk8_270=                    `SPLL_PATH.spll_gen_dclk8_270;
    assign  pll_if.spll_gen_dclk8_315=                    `SPLL_PATH.spll_gen_dclk8_315;
    assign  pll_if.spll_gen_dclk8_45=                     `SPLL_PATH.spll_gen_dclk8_45;
    assign  pll_if.spll_gen_dclk8_90=                     `SPLL_PATH.spll_gen_dclk8_90;
    assign  pll_if.spll_gen_dft_data_out=                 `SPLL_PATH.spll_gen_dft_data_out;
    assign  pll_if.spll_gen_dig_obs_k=                    `SPLL_PATH.spll_gen_dig_obs_k;
    assign  pll_if.spll_gen_dig_obs_kx=                   `SPLL_PATH.spll_gen_dig_obs_kx;
    assign  pll_if.spll_gen_enter_pulse_mode_pllout=      `SPLL_PATH.spll_gen_enter_pulse_mode_pllout;
    assign  pll_if.spll_gen_fall_fbclk_pllout=            `SPLL_PATH.spll_gen_fall_fbclk_pllout;
    assign  pll_if.spll_gen_init_done=                    `SPLL_PATH.spll_gen_init_done;
    assign  pll_if.spll_gen_lowj_clkout_n=                `SPLL_PATH.spll_gen_lowj_clkout_n;
    assign  pll_if.spll_gen_lowj_clkout_p=                `SPLL_PATH.spll_gen_lowj_clkout_p;
    assign  pll_if.spll_gen_obs_trig_k=                   `SPLL_PATH.spll_gen_obs_trig_k;
    assign  pll_if.spll_gen_obs_trig_kx=                  `SPLL_PATH.spll_gen_obs_trig_kx;
    assign  pll_if.spll_gen_pll_charz_h=                  `SPLL_PATH.spll_gen_pll_charz_h;
    assign  pll_if.spll_gen_pll_charz_l=                  `SPLL_PATH.spll_gen_pll_charz_l;
    assign  pll_if.spll_gen_pll_rdy=                      `SPLL_PATH.spll_gen_pll_rdy;
    assign  pll_if.spll_gen_pllout=                       `SPLL_PATH.spll_gen_pllout;
    assign  pll_if.spll_gen_pllout_ack=                   `SPLL_PATH.spll_gen_pllout_ack;
    assign  pll_if.spll_gen_postdiv_ack=                  `SPLL_PATH.spll_gen_postdiv_ack;
    assign  pll_if.spll_gen_pwrok_vddp=                   `SPLL_PATH.spll_gen_pwrok_vddp;
    assign  pll_if.spll_gen_rise_fbclk_dclk4=             `SPLL_PATH.spll_gen_rise_fbclk_dclk4;
    assign  pll_if.spll_gen_rise_fbclk_dclk8=             `SPLL_PATH.spll_gen_rise_fbclk_dclk8;
    assign  pll_if.spll_gen_rise_fbclk_pllout=            `SPLL_PATH.spll_gen_rise_fbclk_pllout;
    assign  pll_if.spll_gen_scan_out=                     `SPLL_PATH.spll_gen_scan_out;
    assign  pll_if.spll_gen_stopmode_gater_dis_pllout=    `SPLL_PATH.spll_gen_stopmode_gater_dis_pllout;
    assign  pll_if.spll_gen_syncbus_out_pllout=           `SPLL_PATH.spll_gen_syncbus_out_pllout;
    assign  pll_if.spll_gen_true_postdiv_pllout=          `SPLL_PATH.spll_gen_true_postdiv_pllout;


`endif
